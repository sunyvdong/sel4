arch arm11

objects {

cnode_client = cnode (2 bits)
cnode_timer = cnode (4 bits)
device_untyped = ut (12 bits, paddr: 0xf8001000) {  }
endpoint = ep
frame = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 122880}])
frame_client_0000 = frame (64k, fill: [{0 65536 CDL_FrameFill_FileData "client" 0}])
frame_client_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 65536}])
frame_client_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 69632}])
frame_client_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 73728}])
frame_client_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 77824}])
frame_client_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 81920}])
frame_client_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 86016}])
frame_client_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 90112}])
frame_client_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 94208}])
frame_client_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 98304}])
frame_client_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 102400}])
frame_client_0011 = frame (4k, fill: [{0 3544 CDL_FrameFill_FileData "client" 106496}])
frame_client_0012 = frame (4k, fill: [{4068 28 CDL_FrameFill_FileData "client" 110564}])
frame_client_0013 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 110592}])
frame_client_0031 = frame (4k, fill: [{0 20 CDL_FrameFill_FileData "client" 184320}])
frame_client_0032 = frame (4k, fill: [])
frame_client_0033 = frame (64k, fill: [])
frame_client_0034 = frame (64k, fill: [])
frame_client_0035 = frame (64k, fill: [])
frame_client_0036 = frame (64k, fill: [])
frame_client_0037 = frame (64k, fill: [])
frame_client_0038 = frame (64k, fill: [])
frame_client_0039 = frame (64k, fill: [])
frame_client_0040 = frame (64k, fill: [])
frame_client_0041 = frame (64k, fill: [])
frame_client_0042 = frame (64k, fill: [])
frame_client_0043 = frame (64k, fill: [])
frame_client_0044 = frame (64k, fill: [])
frame_client_0045 = frame (64k, fill: [])
frame_client_0046 = frame (64k, fill: [])
frame_client_0047 = frame (64k, fill: [])
frame_client_0048 = frame (64k, fill: [])
frame_client_0049 = frame (4k, fill: [])
frame_client_0050 = frame (4k, fill: [])
frame_client_0051 = frame (4k, fill: [])
frame_client_0052 = frame (4k, fill: [])
frame_client_0053 = frame (4k, fill: [])
frame_timer_0000 = frame (64k, fill: [{0 65536 CDL_FrameFill_FileData "timer" 0}])
frame_timer_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 65536}])
frame_timer_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 69632}])
frame_timer_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 73728}])
frame_timer_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 77824}])
frame_timer_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 81920}])
frame_timer_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 86016}])
frame_timer_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 90112}])
frame_timer_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 94208}])
frame_timer_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 98304}])
frame_timer_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 102400}])
frame_timer_0011 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 106496}])
frame_timer_0012 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 110592}])
frame_timer_0013 = frame (4k, fill: [{0 3128 CDL_FrameFill_FileData "timer" 114688}])
frame_timer_0014 = frame (4k, fill: [{4068 28 CDL_FrameFill_FileData "timer" 118756}])
frame_timer_0015 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 118784}])
frame_timer_0034 = frame (4k, fill: [{0 20 CDL_FrameFill_FileData "timer" 196608}])
frame_timer_0035 = frame (4k, fill: [])
frame_timer_0036 = frame (4k, fill: [])
frame_timer_0037 = frame (4k, fill: [])
frame_timer_0038 = frame (4k, fill: [])
frame_timer_0039 = frame (4k, fill: [])
frame_timer_0040 = frame (4k, fill: [])
frame_timer_0041 = frame (4k, fill: [])
frame_timer_0042 = frame (4k, fill: [])
frame_timer_0043 = frame (4k, fill: [])
frame_timer_0044 = frame (4k, fill: [])
frame_timer_0045 = frame (4k, fill: [])
frame_timer_0046 = frame (4k, fill: [])
frame_timer_0047 = frame (4k, fill: [])
frame_timer_0048 = frame (4k, fill: [])
frame_timer_0049 = frame (64k, fill: [])
frame_timer_0050 = frame (64k, fill: [])
frame_timer_0051 = frame (64k, fill: [])
frame_timer_0052 = frame (64k, fill: [])
frame_timer_0053 = frame (64k, fill: [])
frame_timer_0054 = frame (64k, fill: [])
frame_timer_0055 = frame (64k, fill: [])
frame_timer_0056 = frame (64k, fill: [])
frame_timer_0057 = frame (64k, fill: [])
frame_timer_0058 = frame (64k, fill: [])
frame_timer_0059 = frame (64k, fill: [])
frame_timer_0060 = frame (64k, fill: [])
frame_timer_0061 = frame (64k, fill: [])
frame_timer_0062 = frame (64k, fill: [])
frame_timer_0063 = frame (64k, fill: [])
frame_timer_0064 = frame (4k, fill: [])
frame_timer_0065 = frame (4k, fill: [])
frame_timer_0066 = frame (4k, fill: [])
frame_timer_0067 = frame (4k, fill: [])
frame_timer_0068 = frame (4k, fill: [])
frame_timer_0069 = frame (4k, fill: [])
frame_timer_0070 = frame (4k, fill: [])
frame_timer_0071 = frame (4k, fill: [])
ipc_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 180224}])
ipc_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 192512}])
ntfn = notification
pt_client_0000 = pt
pt_client_0046 = pt
pt_timer_0000 = pt
pt_timer_0061 = pt
stack_0_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 114688}])
stack_0_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 126976}])
stack_10_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 155648}])
stack_10_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 167936}])
stack_11_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 159744}])
stack_11_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 172032}])
stack_12_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 163840}])
stack_12_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 176128}])
stack_13_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 167936}])
stack_13_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 180224}])
stack_14_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 172032}])
stack_14_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 184320}])
stack_15_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 176128}])
stack_15_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 188416}])
stack_1_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 118784}])
stack_1_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 131072}])
stack_2_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 122880}])
stack_2_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 135168}])
stack_3_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 126976}])
stack_3_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 139264}])
stack_4_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 131072}])
stack_4_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 143360}])
stack_5_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 135168}])
stack_5_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 147456}])
stack_6_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 139264}])
stack_6_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 151552}])
stack_7_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 143360}])
stack_7_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 155648}])
stack_8_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 147456}])
stack_8_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 159744}])
stack_9_client_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client" 151552}])
stack_9_timer_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "timer" 163840}])
tcb_client = tcb (addr: 0x3d000,ip: 0x10164,sp: 0x2e000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 180232, 1, 0, 0, 32, 76472, 0, 0])
tcb_timer = tcb (addr: 0x40000,ip: 0x10164,sp: 0x31000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 188456, 1, 0, 0, 32, 83424, 0, 0])
vspace_client = pd
vspace_timer = pd
}

caps {
cnode_client {
0x1: endpoint (RWG, badge: 61)
0x2: tcb_client
}
cnode_timer {
0x1: endpoint (RWG)
0x2: ntfn (RWG)
0x3: device_untyped
0x5: cnode_timer (guard: 0, guard_size: 28)
0x6: vspace_timer
0x7: frame (RWX)
0x8: irq_control
0xa: tcb_timer
}
pt_client_0000 {
0x10: frame_client_0000 (RX)
0x20: frame_client_0001 (RX)
0x21: frame_client_0002 (RX)
0x22: frame_client_0003 (RX)
0x23: frame_client_0004 (RX)
0x24: frame_client_0005 (RX)
0x25: frame_client_0006 (RX)
0x26: frame_client_0007 (RX)
0x27: frame_client_0008 (RX)
0x28: frame_client_0009 (RX)
0x29: frame_client_0010 (RX)
0x2a: frame_client_0011 (RX)
0x2b: frame_client_0012 (RW)
0x2c: frame_client_0013 (RW)
0x2d: stack_0_client_obj (RW)
0x2e: stack_1_client_obj (RW)
0x2f: stack_2_client_obj (RW)
0x30: stack_3_client_obj (RW)
0x31: stack_4_client_obj (RW)
0x32: stack_5_client_obj (RW)
0x33: stack_6_client_obj (RW)
0x34: stack_7_client_obj (RW)
0x35: stack_8_client_obj (RW)
0x36: stack_9_client_obj (RW)
0x37: stack_10_client_obj (RW)
0x38: stack_11_client_obj (RW)
0x39: stack_12_client_obj (RW)
0x3a: stack_13_client_obj (RW)
0x3b: stack_14_client_obj (RW)
0x3c: stack_15_client_obj (RW)
0x3d: ipc_client_obj (RW)
0x3e: frame_client_0031 (RW)
0x3f: frame_client_0032 (RW)
0x40: frame_client_0033 (RW)
0x50: frame_client_0034 (RW)
0x60: frame_client_0035 (RW)
0x70: frame_client_0036 (RW)
0x80: frame_client_0037 (RW)
0x90: frame_client_0038 (RW)
0xa0: frame_client_0039 (RW)
0xb0: frame_client_0040 (RW)
0xc0: frame_client_0041 (RW)
0xd0: frame_client_0042 (RW)
0xe0: frame_client_0043 (RW)
0xf0: frame_client_0044 (RW)
}
pt_client_0046 {
0x0: frame_client_0045 (RW)
0x10: frame_client_0046 (RW)
0x20: frame_client_0047 (RW)
0x30: frame_client_0048 (RW)
0x40: frame_client_0049 (RW)
0x41: frame_client_0050 (RW)
0x42: frame_client_0051 (RW)
0x43: frame_client_0052 (RW)
0x44: frame_client_0053 (RW)
}
pt_timer_0000 {
0x10: frame_timer_0000 (RX)
0x20: frame_timer_0001 (RX)
0x21: frame_timer_0002 (RX)
0x22: frame_timer_0003 (RX)
0x23: frame_timer_0004 (RX)
0x24: frame_timer_0005 (RX)
0x25: frame_timer_0006 (RX)
0x26: frame_timer_0007 (RX)
0x27: frame_timer_0008 (RX)
0x28: frame_timer_0009 (RX)
0x29: frame_timer_0010 (RX)
0x2a: frame_timer_0011 (RX)
0x2b: frame_timer_0012 (RX)
0x2c: frame_timer_0013 (RX)
0x2d: frame_timer_0014 (RW)
0x2e: frame_timer_0015 (RW)
0x2f: frame (RWX)
0x30: stack_0_timer_obj (RW)
0x31: stack_1_timer_obj (RW)
0x32: stack_2_timer_obj (RW)
0x33: stack_3_timer_obj (RW)
0x34: stack_4_timer_obj (RW)
0x35: stack_5_timer_obj (RW)
0x36: stack_6_timer_obj (RW)
0x37: stack_7_timer_obj (RW)
0x38: stack_8_timer_obj (RW)
0x39: stack_9_timer_obj (RW)
0x3a: stack_10_timer_obj (RW)
0x3b: stack_11_timer_obj (RW)
0x3c: stack_12_timer_obj (RW)
0x3d: stack_13_timer_obj (RW)
0x3e: stack_14_timer_obj (RW)
0x3f: stack_15_timer_obj (RW)
0x40: ipc_timer_obj (RW)
0x41: frame_timer_0034 (RW)
0x42: frame_timer_0035 (RW)
0x43: frame_timer_0036 (RW)
0x44: frame_timer_0037 (RW)
0x45: frame_timer_0038 (RW)
0x46: frame_timer_0039 (RW)
0x47: frame_timer_0040 (RW)
0x48: frame_timer_0041 (RW)
0x49: frame_timer_0042 (RW)
0x4a: frame_timer_0043 (RW)
0x4b: frame_timer_0044 (RW)
0x4c: frame_timer_0045 (RW)
0x4d: frame_timer_0046 (RW)
0x4e: frame_timer_0047 (RW)
0x4f: frame_timer_0048 (RW)
0x50: frame_timer_0049 (RW)
0x60: frame_timer_0050 (RW)
0x70: frame_timer_0051 (RW)
0x80: frame_timer_0052 (RW)
0x90: frame_timer_0053 (RW)
0xa0: frame_timer_0054 (RW)
0xb0: frame_timer_0055 (RW)
0xc0: frame_timer_0056 (RW)
0xd0: frame_timer_0057 (RW)
0xe0: frame_timer_0058 (RW)
0xf0: frame_timer_0059 (RW)
}
pt_timer_0061 {
0x0: frame_timer_0060 (RW)
0x10: frame_timer_0061 (RW)
0x20: frame_timer_0062 (RW)
0x30: frame_timer_0063 (RW)
0x40: frame_timer_0064 (RW)
0x41: frame_timer_0065 (RW)
0x42: frame_timer_0066 (RW)
0x43: frame_timer_0067 (RW)
0x44: frame_timer_0068 (RW)
0x45: frame_timer_0069 (RW)
0x46: frame_timer_0070 (RW)
0x47: frame_timer_0071 (RW)
}
tcb_client {
cspace: cnode_client (guard: 0, guard_size: 30)
ipc_buffer_slot: ipc_client_obj (RW)
vspace: vspace_client
}
tcb_timer {
cspace: cnode_timer (guard: 0, guard_size: 28)
ipc_buffer_slot: ipc_timer_obj (RW)
vspace: vspace_timer
}
vspace_client {
0x0: pt_client_0000
0x1: pt_client_0046
}
vspace_timer {
0x0: pt_timer_0000
0x1: pt_timer_0061
}
}

irq maps {

}